`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/21/2023 04:15:41 AM
// Design Name: 
// Module Name: tb_crank_cam_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_crank_cam_sim(

    );
    
    
    
    crank_cam_sim_v1_0 crank_cam_sim_v1_0_inst() ;
    
    initial begin
    #100 finish;
    end
endmodule
